module ring(input )